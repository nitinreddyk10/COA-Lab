module not_v (input a, output out);
    not (out, a);
endmodule
